-- TestSystem
--
-- Combine the ByteMachine together with a proper ROM
-- and set up output ports for the test program to produce some signals.AD/STORE operations)

library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

use work.ByteMachine_pkg.all;

entity TestSystem is	
	port (
		clk: in std_logic;		
		reset: in std_logic;  -- active low!
		
		-- ouput ports
		port0 : out unsigned(7 downto 0);
		
		-- test output
		test_pc : out unsigned(15 downto 0);
		test_sp : out unsigned(7 downto 0);
		test_r : out unsigned(7 downto 0);
		test_fetchb : out std_logic
	);
		
end entity;

architecture rtl of TestSystem is

	component ByteMachine
	generic ( 
		 numinputports:integer;
		 numoutputports:integer;
		 code:bytemachinecode
	 );
	port (
		clk: in std_logic;		
		reset: in std_logic;
				
		-- ports
		input : in bytemachineports(0 to numinputports-1);
		output : out bytemachineports(0 to numoutputports-1);
				
		-- test output
		test_pc : out unsigned(15 downto 0);
		test_sp : out unsigned(7 downto 0);
		test_r : out unsigned(7 downto 0);
		test_fetchb : out std_logic
	);
	end component;		
	
   constant code : bytemachinecode := ( 
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,
16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,
16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,
16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#13#,16#10#,16#00#,16#DE#,16#20#,16#12#,16#0E#,
16#10#,16#00#,16#E0#,16#1D#,16#12#,16#00#,16#D2#,16#20#,16#18#,16#10#,16#00#,16#DF#,16#20#,16#10#,16#12#,16#00#,
16#D9#,16#20#,16#17#,16#12#,16#00#,16#DC#,16#20#,16#E1#,16#1C#,16#1D#,16#04#,16#11#,16#06#,16#12#,16#07#,16#19#,
16#07#,16#10#,16#02#,16#18#,16#06#,16#11#,16#06#,16#14#,16#06#,16#10#,16#02#,16#11#,16#06#,16#10#,16#02#,16#1C#,
16#06#,16#15#,16#12#,16#00#,16#D2#,16#20#,16#1C#,16#19#,16#06#,16#14#,16#07#,16#14#,16#07#,16#1C#,16#06#,16#15#,
16#06#,16#10#,16#02#,16#1C#,16#06#,16#11#,16#06#,16#1D#,16#06#,16#12#,16#06#,16#1C#,16#02#,16#10#,16#02#,16#15#,
16#12#,16#00#,16#D2#,16#20#,16#1C#,16#18#,16#04#,16#19#,16#06#,16#13#,16#07#,16#10#,16#02#,16#16#,16#06#,16#1C#,
16#06#,16#15#,16#06#,16#15#,16#06#,16#13#,16#06#,16#15#,16#06#,16#10#,16#02#,16#17#,16#07#,16#15#,16#12#,16#00#,
16#D2#,16#20#,16#1C#,16#11#,16#06#,16#13#,16#07#,16#10#,16#02#,16#17#,16#07#,16#18#,16#06#,16#19#,16#06#,16#14#,
16#07#,16#15#,16#06#,16#10#,16#02#,16#11#,16#06#,16#13#,16#07#,16#10#,16#02#,16#15#,16#12#,16#00#,16#D2#,16#20#,
16#1C#,16#13#,16#07#,16#1E#,16#06#,16#1F#,16#06#,16#17#,16#07#,16#1C#,16#02#,16#10#,16#02#,16#11#,16#04#,16#1E#,
16#06#,16#14#,16#06#,16#10#,16#02#,16#15#,16#06#,16#16#,16#07#,16#15#,16#12#,16#00#,16#D2#,16#20#,16#1C#,16#15#,
16#06#,16#12#,16#07#,16#19#,16#07#,16#17#,16#07#,16#18#,16#06#,16#15#,16#06#,16#12#,16#07#,16#15#,16#06#,16#10#,
16#02#,16#14#,16#07#,16#18#,16#06#,16#11#,16#06#,16#15#,16#12#,16#00#,16#D2#,16#20#,16#1C#,16#14#,16#07#,16#10#,
16#02#,16#1D#,16#04#,16#11#,16#06#,16#12#,16#07#,16#19#,16#07#,16#10#,16#02#,16#17#,16#07#,16#15#,16#06#,16#1E#,
16#06#,16#14#,16#07#,16#1C#,16#02#,16#15#,16#12#,16#00#,16#D2#,16#20#,16#1C#,16#10#,16#02#,16#14#,16#05#,16#18#,
16#06#,16#15#,16#06#,16#10#,16#02#,16#1C#,16#06#,16#11#,16#06#,16#1D#,16#06#,16#12#,16#06#,16#10#,16#02#,16#17#,
16#07#,16#11#,16#06#,16#15#,16#12#,16#00#,16#D2#,16#20#,16#1C#,16#13#,16#07#,16#10#,16#02#,16#13#,16#07#,16#15#,
16#07#,16#12#,16#07#,16#15#,16#06#,16#10#,16#02#,16#14#,16#07#,16#1F#,16#06#,16#10#,16#02#,16#17#,16#06#,16#1F#,
16#06#,16#15#,16#12#,16#00#,16#D2#,16#20#,16#11#,16#1E#,16#02#,16#18#,16#07#,16#18#,16#07#,16#18#,16#07#,16#18#,
16#07#,16#18#,16#07#,16#18#,16#07#,16#18#,16#07#,16#18#,16#07#,16#18#,16#07#,16#18#,16#07#,16#18#,16#07#,16#15#,
16#12#,16#00#,16#D2#,16#20#,16#E1#,16#3D#,16#4F#,16#1A#,16#12#,16#00#,16#D7#,16#20#,16#EE#,16#11#,16#00#,16#13#,
16#02#,16#15#,16#04#,16#17#,16#06#,16#10#,16#15#,16#18#,16#00#,16#D7#,16#20#,16#19#,16#08#,16#1B#,16#0A#,16#1D#,
16#0C#,16#1F#,16#0E#,16#14#,16#15#,16#18#,16#00#,16#D7#,16#20#,16#1E#,16#0F#,16#1C#,16#0D#,16#1A#,16#0B#,16#18#,
16#09#,16#18#,16#15#,16#18#,16#00#,16#D7#,16#20#,16#16#,16#07#,16#14#,16#05#,16#12#,16#03#,16#10#,16#01#,16#1C#,
16#15#,16#18#,16#00#,16#D7#,16#20#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#11#,16#05#,16#15#,
16#18#,16#00#,16#D7#,16#20#,16#10#,16#10#,16#05#,16#70#,16#20#,16#E1#,16#42#,16#C0#,16#E3#,16#43#,16#60#,16#11#,
16#15#,16#12#,16#00#,16#DE#,16#20#,16#43#,16#11#,16#21#,16#53#,16#42#,16#11#,16#22#,16#52#,16#1E#,16#0F#,16#AB#,
16#10#,16#08#,16#10#,16#15#,16#12#,16#00#,16#DE#,16#20#,16#10#,16#05#,16#60#,16#18#,16#03#,16#25#,16#B9#,16#10#,
16#10#,16#15#,16#12#,16#00#,16#DE#,16#20#,16#1F#,16#0F#,16#A0#,16#11#,16#05#,16#18#,16#04#,16#1D#,16#18#,16#00#,
16#D7#,16#20#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#10#,16#00#,16#1C#,16#04#,16#15#,16#18#,16#00#,16#D7#,
16#20#,16#10#,16#13#,16#00#,16#D2#,16#20#,16#E1#,16#10#,16#1B#,16#19#,16#00#,16#D7#,16#20#,16#14#,16#1B#,16#19#,
16#00#,16#D7#,16#20#,16#18#,16#1B#,16#19#,16#00#,16#D7#,16#20#,16#1C#,16#1B#,16#19#,16#00#,16#D7#,16#20#,16#14#,
16#19#,16#00#,16#D7#,16#20#,16#E1#,16#42#,16#C2#,16#11#,16#00#,16#A5#,16#18#,16#00#,16#10#,16#00#,16#10#,16#00#,
16#10#,16#00#,16#33#,16#11#,16#05#,16#15#,16#18#,16#00#,16#DF#,16#20#,16#20#,16#20#,16#20#,16#20#,16#43#,16#10#,
16#05#,16#60#,16#10#,16#01#,16#21#,16#70#,16#20#,16#10#,16#05#,16#60#,16#11#,16#21#,16#40#,16#10#,16#05#,16#70#,
16#20#,16#10#,16#04#,16#25#,16#C9#,16#10#,16#13#,16#00#,16#D2#,16#20#,16#10#,16#10#,16#05#,16#70#,16#20#,16#E3#,
16#10#,16#15#,16#05#,16#1D#,16#18#,16#00#,16#D7#,16#20#,16#14#,16#19#,16#05#,16#1D#,16#18#,16#00#,16#D7#,16#20#,
16#18#,16#1D#,16#05#,16#1D#,16#18#,16#00#,16#D7#,16#20#,16#1C#,16#11#,16#06#,16#1D#,16#18#,16#00#,16#D7#,16#20#,
16#18#,16#07#,16#14#,16#0A#,16#1A#,16#06#,16#17#,16#0D#,16#17#,16#10#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#16#,
16#05#,16#17#,16#0B#,16#17#,16#0C#,16#18#,16#0E#,16#1C#,16#11#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#1B#,16#0D#,
16#10#,16#07#,16#10#,16#02#,16#14#,16#02#,16#11#,16#01#,16#12#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#1E#,16#0E#,
16#1E#,16#0C#,16#1D#,16#0B#,16#11#,16#0C#,16#16#,16#01#,16#13#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#1F#,16#0A#,
16#1F#,16#00#,16#1C#,16#07#,16#15#,16#0F#,16#17#,16#14#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#1A#,16#02#,16#16#,
16#0C#,16#17#,16#08#,16#17#,16#04#,16#1C#,16#15#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#13#,16#01#,16#16#,16#04#,
16#10#,16#03#,16#18#,16#0A#,16#11#,16#01#,16#16#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#11#,16#00#,16#15#,16#09#,
16#16#,16#04#,16#1D#,16#0F#,16#16#,16#01#,16#17#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#18#,16#0D#,16#18#,16#09#,
16#10#,16#08#,16#19#,16#06#,16#17#,16#18#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#1F#,16#0A#,16#17#,16#0F#,16#14#,
16#04#,16#1B#,16#08#,16#1C#,16#19#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#11#,16#0B#,16#1B#,16#05#,16#1F#,16#0F#,
16#1F#,16#0F#,16#11#,16#01#,16#1A#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#1E#,16#0B#,16#17#,16#0D#,16#1C#,16#05#,
16#19#,16#08#,16#16#,16#01#,16#1B#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#12#,16#02#,16#11#,16#01#,16#10#,16#09#,
16#1B#,16#06#,16#17#,16#1C#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#13#,16#09#,16#11#,16#07#,16#18#,16#09#,16#1D#,
16#0F#,16#1C#,16#1D#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#1E#,16#08#,16#13#,16#04#,16#19#,16#07#,16#16#,16#0A#,
16#11#,16#01#,16#1E#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#11#,16#02#,16#18#,16#00#,16#14#,16#0B#,16#19#,16#04#,
16#16#,16#01#,16#1F#,16#19#,16#17#,16#00#,16#D3#,16#20#,16#12#,16#06#,16#15#,16#02#,16#1E#,16#01#,16#16#,16#0F#,
16#15#,16#11#,16#16#,16#17#,16#00#,16#D6#,16#20#,16#10#,16#04#,16#13#,16#0B#,16#10#,16#04#,16#10#,16#0C#,16#19#,
16#16#,16#16#,16#17#,16#00#,16#D6#,16#20#,16#11#,16#05#,16#1A#,16#05#,16#1E#,16#05#,16#16#,16#02#,16#1E#,16#1B#,
16#16#,16#17#,16#00#,16#D6#,16#20#,16#1A#,16#0A#,16#17#,16#0C#,16#16#,16#0B#,16#19#,16#0E#,16#14#,16#01#,16#10#,
16#16#,16#17#,16#00#,16#D6#,16#20#,16#1D#,16#05#,16#10#,16#01#,16#1F#,16#02#,16#16#,16#0D#,16#15#,16#15#,16#16#,
16#17#,16#00#,16#D6#,16#20#,16#13#,16#05#,16#14#,16#01#,16#14#,16#04#,16#12#,16#00#,16#19#,16#1A#,16#16#,16#17#,
16#00#,16#D6#,16#20#,16#11#,16#08#,16#16#,16#0E#,16#11#,16#0A#,16#18#,16#0D#,16#1E#,16#1F#,16#16#,16#17#,16#00#,
16#D6#,16#20#,16#18#,16#0C#,16#1B#,16#0F#,16#13#,16#0D#,16#17#,16#0E#,16#14#,16#01#,16#14#,16#16#,16#17#,16#00#,
16#D6#,16#20#,16#16#,16#0E#,16#1D#,16#0C#,16#11#,16#0E#,16#11#,16#02#,16#15#,16#19#,16#16#,16#17#,16#00#,16#D6#,
16#20#,16#16#,16#0D#,16#17#,16#00#,16#17#,16#03#,16#13#,16#0C#,16#19#,16#1E#,16#16#,16#17#,16#00#,16#D6#,16#20#,
16#17#,16#08#,16#1D#,16#00#,16#15#,16#0D#,16#14#,16#0F#,16#1E#,16#13#,16#16#,16#17#,16#00#,16#D6#,16#20#,16#1D#,
16#0E#,16#14#,16#01#,16#1A#,16#05#,16#15#,16#04#,16#14#,16#01#,16#18#,16#16#,16#17#,16#00#,16#D6#,16#20#,16#15#,
16#00#,16#19#,16#0E#,16#13#,16#0E#,16#19#,16#0A#,16#15#,16#1D#,16#16#,16#17#,16#00#,16#D6#,16#20#,16#18#,16#0F#,
16#13#,16#0A#,16#1F#,16#0E#,16#1C#,16#0F#,16#19#,16#12#,16#16#,16#17#,16#00#,16#D6#,16#20#,16#19#,16#0D#,16#12#,
16#00#,16#1F#,16#06#,16#17#,16#06#,16#1E#,16#17#,16#16#,16#17#,16#00#,16#D6#,16#20#,16#1A#,16#08#,16#1C#,16#04#,
16#1A#,16#02#,16#1D#,16#08#,16#14#,16#01#,16#1C#,16#16#,16#17#,16#00#,16#D6#,16#20#,16#12#,16#04#,16#19#,16#03#,
16#1A#,16#0F#,16#1F#,16#0F#,16#14#,16#15#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#11#,16#08#,16#16#,16#0F#,16#11#,
16#07#,16#17#,16#08#,16#1B#,16#18#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#12#,16#02#,16#11#,16#06#,16#1D#,16#09#,
16#1D#,16#06#,16#10#,16#01#,16#1B#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#1C#,16#00#,16#18#,16#03#,16#15#,16#0E#,
16#1D#,16#0F#,16#17#,16#01#,16#1E#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#14#,16#04#,16#1A#,16#0E#,16#1E#,16#0B#,
16#14#,16#0A#,16#14#,16#11#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#19#,16#0A#,16#1F#,16#0C#,16#1E#,16#0D#,16#1B#,
16#04#,16#1B#,16#14#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#10#,16#06#,16#1B#,16#04#,16#1B#,16#0B#,16#16#,16#0F#,
16#10#,16#01#,16#17#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#10#,16#07#,16#1C#,16#0B#,16#1F#,16#0B#,16#1E#,16#0B#,
16#17#,16#01#,16#1A#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#16#,16#0C#,16#1E#,16#07#,16#1B#,16#09#,16#18#,16#02#,
16#14#,16#1D#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#1A#,16#0F#,16#17#,16#02#,16#11#,16#0A#,16#1A#,16#0E#,16#1B#,
16#10#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#15#,16#08#,16#10#,16#03#,16#1F#,16#0E#,16#14#,16#0D#,16#10#,16#01#,
16#13#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#15#,16#00#,16#1D#,16#01#,16#18#,16#08#,16#14#,16#00#,16#17#,16#01#,
16#16#,16#13#,16#17#,16#00#,16#D9#,16#20#,16#19#,16#03#,16#10#,16#0D#,16#14#,16#0D#,16#19#,16#0D#,16#14#,16#19#,
16#13#,16#17#,16#00#,16#D9#,16#20#,16#15#,16#0E#,16#19#,16#09#,16#1B#,16#0D#,16#16#,16#0E#,16#1B#,16#1C#,16#13#,
16#17#,16#00#,16#D9#,16#20#,16#18#,16#0F#,16#1C#,16#07#,16#12#,16#0A#,16#1F#,16#01#,16#10#,16#01#,16#1F#,16#13#,
16#17#,16#00#,16#D9#,16#20#,16#15#,16#06#,16#16#,16#05#,16#1C#,16#0A#,16#14#,16#0C#,16#17#,16#01#,16#12#,16#13#,
16#17#,16#00#,16#D9#,16#20#,16#14#,16#04#,16#12#,16#02#,16#19#,16#02#,16#14#,16#0F#,16#16#,16#10#,16#17#,16#17#,
16#00#,16#DB#,16#20#,16#17#,16#09#,16#1F#,16#0F#,16#1A#,16#02#,16#13#,16#04#,16#1A#,16#17#,16#17#,16#17#,16#00#,
16#DB#,16#20#,16#17#,16#0A#,16#13#,16#02#,16#14#,16#09#,16#1B#,16#0A#,16#1F#,16#1E#,16#17#,16#17#,16#00#,16#DB#,
16#20#,16#19#,16#03#,16#10#,16#0A#,16#13#,16#09#,16#1C#,16#0F#,16#15#,16#01#,16#15#,16#17#,16#17#,16#00#,16#DB#,
16#20#,16#13#,16#0C#,16#19#,16#05#,16#1B#,16#05#,16#15#,16#06#,16#16#,16#1C#,16#17#,16#17#,16#00#,16#DB#,16#20#,
16#12#,16#09#,16#1C#,16#0C#,16#1C#,16#00#,16#1F#,16#08#,16#1A#,16#13#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#1D#,
16#07#,16#14#,16#0F#,16#1F#,16#0E#,16#1F#,16#0F#,16#1F#,16#1A#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#11#,16#0D#,
16#1D#,16#05#,16#14#,16#08#,16#15#,16#08#,16#15#,16#01#,16#11#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#1F#,16#04#,
16#1E#,16#07#,16#18#,16#0A#,16#1F#,16#06#,16#16#,16#18#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#10#,16#0E#,16#16#,
16#0E#,16#1C#,16#02#,16#1E#,16#0F#,16#1A#,16#1F#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#14#,16#01#,16#13#,16#04#,
16#11#,16#00#,16#13#,16#0A#,16#1F#,16#16#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#11#,16#0A#,16#11#,16#01#,16#18#,
16#00#,16#1E#,16#04#,16#15#,16#01#,16#1D#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#12#,16#08#,16#1E#,16#07#,16#13#,
16#05#,16#17#,16#0F#,16#16#,16#14#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#15#,16#03#,16#12#,16#0F#,16#1A#,16#03#,
16#1D#,16#0B#,16#1A#,16#1B#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#1B#,16#0B#,16#12#,16#0D#,16#17#,16#0D#,16#1A#,
16#02#,16#1F#,16#12#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#11#,16#09#,16#13#,16#0D#,16#16#,16#08#,16#1B#,16#0E#,
16#15#,16#01#,16#19#,16#17#,16#17#,16#00#,16#DB#,16#20#,16#15#,16#05#,16#10#,16#15#,16#18#,16#00#,16#DF#,16#20#,
16#19#,16#05#,16#14#,16#15#,16#18#,16#00#,16#DF#,16#20#,16#1D#,16#05#,16#18#,16#15#,16#18#,16#00#,16#DF#,16#20#,
16#11#,16#06#,16#1C#,16#15#,16#18#,16#00#,16#DF#,16#20#,16#E1#,16#1D#,16#05#,16#19#,16#06#,16#1D#,16#18#,16#00#,
16#D7#,16#20#,16#11#,16#06#,16#19#,16#06#,16#14#,16#18#,16#00#,16#DD#,16#20#,16#19#,16#05#,16#19#,16#06#,16#12#,
16#18#,16#00#,16#D9#,16#20#,16#11#,16#06#,16#19#,16#06#,16#14#,16#18#,16#00#,16#DD#,16#20#,16#37#,16#44#,16#44#,
16#1F#,16#18#,16#00#,16#D1#,16#20#,16#E7#,16#19#,16#05#,16#19#,16#06#,16#1D#,16#18#,16#00#,16#D7#,16#20#,16#1D#,
16#05#,16#19#,16#06#,16#14#,16#18#,16#00#,16#DD#,16#20#,16#11#,16#06#,16#19#,16#06#,16#12#,16#18#,16#00#,16#D9#,
16#20#,16#1D#,16#05#,16#19#,16#06#,16#14#,16#18#,16#00#,16#DD#,16#20#,16#37#,16#44#,16#44#,16#1F#,16#18#,16#00#,
16#D1#,16#20#,16#E7#,16#19#,16#05#,16#19#,16#06#,16#1D#,16#18#,16#00#,16#D7#,16#20#,16#1D#,16#05#,16#19#,16#06#,
16#14#,16#18#,16#00#,16#DD#,16#20#,16#11#,16#06#,16#19#,16#06#,16#14#,16#18#,16#00#,16#DD#,16#20#,16#37#,16#44#,
16#44#,16#1F#,16#18#,16#00#,16#D1#,16#20#,16#E7#,16#1F#,16#0F#,16#1F#,16#0F#,16#1F#,16#0F#,16#1F#,16#0F#,16#33#,
16#19#,16#06#,16#1D#,16#18#,16#00#,16#D7#,16#20#,16#20#,16#20#,16#20#,16#20#,16#11#,16#06#,16#19#,16#06#,16#14#,
16#18#,16#00#,16#DD#,16#20#,16#19#,16#05#,16#19#,16#06#,16#13#,16#18#,16#00#,16#DB#,16#20#,16#1D#,16#05#,16#19#,
16#06#,16#14#,16#18#,16#00#,16#DD#,16#20#,16#37#,16#44#,16#44#,16#1F#,16#18#,16#00#,16#D1#,16#20#,16#E7#,16#15#,
16#05#,16#1B#,16#19#,16#00#,16#D7#,16#20#,16#19#,16#05#,16#1B#,16#19#,16#00#,16#D7#,16#20#,16#1D#,16#05#,16#1B#,
16#19#,16#00#,16#D7#,16#20#,16#11#,16#06#,16#1B#,16#19#,16#00#,16#D7#,16#20#,16#19#,16#06#,16#1B#,16#19#,16#00#,
16#D7#,16#20#,16#15#,16#06#,16#1B#,16#19#,16#00#,16#D7#,16#20#,16#14#,16#19#,16#00#,16#D7#,16#20#,16#E1#,16#44#,
16#15#,16#06#,16#1D#,16#18#,16#00#,16#D7#,16#20#,16#15#,16#05#,16#19#,16#06#,16#15#,16#18#,16#00#,16#DF#,16#20#,
16#15#,16#06#,16#19#,16#06#,16#15#,16#18#,16#00#,16#DF#,16#20#,16#10#,16#01#,16#43#,16#10#,16#28#,16#10#,16#28#,
16#21#,16#19#,16#06#,16#15#,16#18#,16#00#,16#DF#,16#20#,16#43#,16#19#,16#06#,16#19#,16#19#,16#00#,16#D4#,16#20#,
16#11#,16#06#,16#15#,16#05#,16#1D#,16#18#,16#00#,16#D7#,16#20#,16#1D#,16#05#,16#11#,16#06#,16#1D#,16#18#,16#00#,
16#D7#,16#20#,16#19#,16#05#,16#1D#,16#05#,16#1D#,16#18#,16#00#,16#D7#,16#20#,16#19#,16#06#,16#19#,16#05#,16#15#,
16#18#,16#00#,16#DF#,16#20#,16#E4#,16#36#,16#43#,16#1D#,16#18#,16#00#,16#D7#,16#20#,16#E6#,16#43#,16#60#,16#43#,
16#70#,16#20#,16#43#,16#61#,16#43#,16#71#,16#20#,16#43#,16#62#,16#43#,16#72#,16#20#,16#43#,16#63#,16#43#,16#73#,
16#20#,16#E3#,16#43#,16#60#,16#43#,16#60#,16#23#,16#43#,16#70#,16#20#,16#43#,16#61#,16#43#,16#61#,16#23#,16#43#,
16#71#,16#20#,16#43#,16#62#,16#43#,16#62#,16#23#,16#43#,16#72#,16#20#,16#43#,16#63#,16#43#,16#63#,16#23#,16#43#,
16#73#,16#20#,16#E3#,16#43#,16#60#,16#43#,16#60#,16#24#,16#43#,16#70#,16#20#,16#43#,16#61#,16#43#,16#61#,16#24#,
16#43#,16#71#,16#20#,16#43#,16#62#,16#43#,16#62#,16#24#,16#43#,16#72#,16#20#,16#43#,16#63#,16#43#,16#63#,16#24#,
16#43#,16#73#,16#20#,16#E3#,16#43#,16#60#,16#43#,16#60#,16#25#,16#43#,16#70#,16#20#,16#43#,16#61#,16#43#,16#61#,
16#25#,16#43#,16#71#,16#20#,16#43#,16#62#,16#43#,16#62#,16#25#,16#43#,16#72#,16#20#,16#43#,16#63#,16#43#,16#63#,
16#25#,16#43#,16#73#,16#20#,16#E3#,16#10#,16#44#,16#60#,16#44#,16#60#,16#18#,16#19#,16#00#,16#D2#,16#20#,16#44#,
16#70#,16#20#,16#44#,16#61#,16#44#,16#61#,16#18#,16#19#,16#00#,16#D2#,16#20#,16#44#,16#71#,16#20#,16#44#,16#62#,
16#44#,16#62#,16#18#,16#19#,16#00#,16#D2#,16#20#,16#44#,16#72#,16#20#,16#44#,16#63#,16#44#,16#63#,16#18#,16#19#,
16#00#,16#D2#,16#20#,16#44#,16#73#,16#20#,16#20#,16#E3#,16#43#,16#43#,16#1F#,16#0F#,16#25#,16#27#,16#B8#,16#43#,
16#43#,16#21#,16#45#,16#21#,16#53#,16#11#,16#54#,16#E2#,16#43#,16#43#,16#21#,16#53#,16#44#,16#C0#,16#E2#,16#11#,
16#44#,16#21#,16#53#,16#43#,16#C0#,16#E2#,16#10#,16#54#,16#E2#,16#43#,16#C0#,16#E3#,16#42#,16#63#,16#40#,16#44#,
16#62#,16#28#,16#44#,16#73#,16#20#,16#43#,16#62#,16#44#,16#61#,16#28#,16#44#,16#72#,16#20#,16#43#,16#61#,16#44#,
16#60#,16#28#,16#44#,16#71#,16#20#,16#43#,16#60#,16#41#,16#28#,16#44#,16#70#,16#20#,16#20#,16#43#,16#11#,16#22#,
16#53#,16#1D#,16#0F#,16#A6#,16#1A#,16#12#,16#19#,16#00#,16#DC#,16#20#,16#E1#,16#42#,16#60#,16#18#,16#19#,16#00#,
16#D9#,16#20#,16#42#,16#61#,16#18#,16#19#,16#00#,16#D9#,16#20#,16#42#,16#62#,16#18#,16#19#,16#00#,16#D9#,16#20#,
16#42#,16#63#,16#18#,16#19#,16#00#,16#D9#,16#20#,16#E2#,16#42#,16#10#,16#29#,16#10#,16#29#,16#10#,16#29#,16#10#,
16#29#,16#1F#,16#19#,16#00#,16#DA#,16#20#,16#42#,16#1F#,16#23#,16#1F#,16#19#,16#00#,16#DA#,16#20#,16#E2#,16#42#,
16#10#,16#03#,16#21#,16#1A#,16#03#,16#41#,16#41#,16#26#,16#50#,16#C1#,16#17#,16#21#,16#12#,16#19#,16#00#,16#DC#,
16#20#,16#E2#,16#42#,16#9F#,16#E2#
	);
begin		
	bm: ByteMachine   
	        generic map(1,1,code) 
	        port map (clk=>clk,
			            reset=>reset, 
							input(0)=>"00000000",
							output(0)=>port0,
	                  test_pc=>test_pc,
							test_sp=>test_sp,
							test_r=>test_r,
							test_fetchb=>test_fetchb);
	
end rtl;


