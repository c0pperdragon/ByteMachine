library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

package Globals is   
	
						
end Globals;

package body Globals is
   -- subprogram bodies here
end Globals;
