-- ByteMachine

library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

package ByteMachine_pkg is
	type bytemachinecode is array(natural range <>) of integer range 0 to 255;
   type bytemachineports is array(natural range <>) of unsigned(7 downto 0);
end package;


library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.ByteMachine_pkg.all;


entity ByteMachine is	
	generic ( 
		 numinputports:integer;
		 numoutputports:integer;
		 code:bytemachinecode
	 );
	port (
		clk: in std_logic;		
		reset: in std_logic;
				
		-- ports
		input : in bytemachineports(0 to numinputports-1);
		output : out bytemachineports(0 to numoutputports-1);
				
		-- test output
		test_pc : out unsigned(15 downto 0);
		test_sp : out unsigned(7 downto 0);
		test_r : out unsigned(7 downto 0);
		test_fetchb : out std_logic
	);
end entity;


architecture rtl of ByteMachine is

	component ByteRAM
	port (
		clk: in std_logic;		
		readaddress : in unsigned(7 downto 0);	
		readdata: out unsigned(7 downto 0);	
		writeaddress : in unsigned(7 downto 0);	
		writedata: in unsigned(7 downto 0);	
		we: in std_logic  );
	end component;		

	component ByteROM
	generic ( 
		 code: bytemachinecode
	);
	PORT
	(
		clock		: IN STD_LOGIC  := '1';
		address		: IN unsigned (15 DOWNTO 0);
		q		    : OUT unsigned (7 DOWNTO 0)
	);
	end component;		
	
	component ByteALU
	port (
		OP: in unsigned (3 downto 0);
		A: in unsigned (7 downto 0);	
		B: in unsigned (7 downto 0);	
		X: out unsigned(7 downto 0)
	);	
	end component;	
		
	-- signals to communicate with the components 
	signal readaddress : unsigned(7 downto 0);	
	signal readdata: unsigned(7 downto 0);	
	signal writeaddress : unsigned(7 downto 0);	
	signal writedata: unsigned(7 downto 0);	
	signal we : std_logic;	

	signal romaddress: unsigned(15 downto 0);
	signal romdata: unsigned(7 downto 0);

	signal aluop : unsigned(3 downto 0);
	signal alua : unsigned(7 downto 0);
	signal alub : unsigned(7 downto 0);
	signal alux : unsigned(7 downto 0);
	 
begin		
	ram: ByteRAM 	
			port map (clk,readaddress,readdata,writeaddress,writedata,we);
	rom: ByteROM 
	      generic map(code) 
	      port map (clk, romaddress, romdata);
	alu: ByteALU
			port map (aluop,alua,alub,alux);
	
	------------------------------- CPU process ------------------
	process (clk,reset,romdata,readdata,alux,input)			
	-- registers
	variable PC : unsigned (15 downto 0) := "0000000000000000";	
	variable SP : unsigned(7 downto 0) := "11111111";
	variable R : unsigned(7 downto 0) := "00000000";
	variable FETCHB : std_logic := '0';
	variable O : bytemachineports(0 to numoutputports-1) := (others => "11111111");
	
	-- temporary variables
	variable A : unsigned(7 downto 0);
	variable B : unsigned(7 downto 0);
	variable opcode : integer range 0 to 15;
	variable x : integer range 0 to 15;
	variable tmp12 : unsigned(11 downto 0);
	variable tmp16 : unsigned(15 downto 0);
	variable pcnew : unsigned (15 downto 0);
	
	-- flags generated by the decoding stage ---
	variable R_NEW : unsigned(7 downto 0);
	variable FETCHB_NEW : std_logic;
	type pcchange_t is (pcinc,pcbranch,pcnear,pcfar);
	variable PCCHANGE : pcchange_t;
	type spchange_t is (spnop,spinc,spdec,spdecx);
	variable SPCHANGE : spchange_t;
	variable WRITEOUT : boolean;
	
	begin			
		----------- asynchronious logic ---------------
		-- decide from where the operands must be taken
		if FETCHB='1' then 
			A := R;
			B := readdata; 
		else
			A := readdata;
			B := R; 	
		end if;
		
		-- feed correct operands into alu --
		aluop <= romdata(3 downto 0);
		alua <= A;
		alub <= B;
		
		-- default flags for execution stage ----
		R_NEW := B;
		FETCHB_NEW := '0';
		PCCHANGE := pcinc;
		SPCHANGE := spnop; 
		WRITEOUT := false;

		-- default values for ram interface --
		readaddress <= SP-1; -- "00000000"; // unsigned(7 downto 0);	
		writeaddress <= SP; -- 00000000"; // : unsigned(7 downto 0);	
		writedata <= B; --: unsigned(7 downto 0);	
		we <= '0'; -- : std_logic;	

		-- decode instruction (also setting some outgoing signals) --
		opcode := to_integer(romdata(7 downto 4));
		x := to_integer(romdata(3 downto 0));
		case opcode is
		when 0 =>    -- EXT x
			R_NEW := (romdata(3 downto 0) or B(7 downto 4)) & B(3 downto 0);
			readaddress <= SP-1;
			SPCHANGE := spnop;
		when 1 =>    -- DAT x
			R_NEW := "0000" & romdata(3 downto 0);
			writeaddress <= SP;
			writedata <= B;
			we <='1';
			readaddress <= SP;
			SPCHANGE := spinc;
	   when 2 => -- OP x
			R_NEW := alux;
			readaddress <= SP-2;
			SPCHANGE := spdec;
		when 3 => -- ADR x
			R_NEW := SP - x;
			writeaddress <= SP;
			writedata <= B;
			we <='1';
			readaddress <= SP;
			SPCHANGE := spinc;
		when 4 => -- GET x
			R_NEW := B;
			FETCHB_NEW := '1';
			writeaddress <= SP;
			writedata <= B;
			we <='1';
			readaddress <= SP-x;
			SPCHANGE := spinc;
		when 5 => -- SET x
			R_NEW := A;
			if x=0 then
				R_NEW := B;
			end if;
			writeaddress <= SP - 1 - x;
			writedata <= B;
			we <='1';
			readaddress <= SP-2;
			SPCHANGE := spdec;
		when 6 => -- LOD x
			R_NEW := A;
			FETCHB_NEW := '1';
			writeaddress <= SP;
			writedata <= B;
			we <='1';
			readaddress <= B + x;			
			SPCHANGE := spnop;		
		when 7 => -- STO x
			R_NEW := A;
			writeaddress <= B + x;
			writedata <= A;
			we <= '1';
			readaddress <= SP-2;
			SPCHANGE := spdec;			
		when 8 => -- IN x
			R_NEW := input(x);
			writeaddress <= SP;
			writedata <= B;
			we <='1';
			readaddress <= SP;
			SPCHANGE := spinc;		
		when 9 => -- OUT x
			WRITEOUT := true;
			R_NEW := A;
			readaddress <= SP-2;
			SPCHANGE := spdec;
		when 10 => -- JMP x
			R_NEW := A;
			readaddress <= SP-2;
			SPCHANGE := spdec;
			PCCHANGE := pcnear;
		when 11 => -- JZ x
			R_NEW := A;
			readaddress <= SP-2; 
			SPCHANGE := spdec;
			if B="00000000" then 
				PCCHANGE := pcbranch;
			end if;
		when 12 => -- JNZ x
			R_NEW := A;
			readaddress <= SP-2; 
			SPCHANGE := spdec;
			if B/="00000000" then 
				PCCHANGE := pcbranch;
			end if;
		when 13 => -- JSR x
			tmp16 := PC+1;
			R_NEW := tmp16(15 downto 8);
			readaddress <= SP-1;
			writeaddress <= SP - 1;
			writedata <= tmp16(7 downto 0);
			we <= '1';
			SPCHANGE := spnop;
			PCCHANGE := pcfar; 
		when 14 => -- RET x
			R_NEW := B;
			readaddress <= SP-x-1; 
			SPCHANGE := spdecx;
			PCCHANGE := pcfar; 
		when 15 => -- reserved
		end case;
		
		-------- determine next instruction address --------
		case PCCHANGE is
		when pcinc => pcnew := PC+1;
		when pcbranch => pcnew := PC + 2 + x;
		when pcnear =>
			tmp12 := B & to_unsigned(x,4); 
			pcnew:= PC + (tmp12(11 downto 11) & tmp12(11) & tmp12(11) & tmp12(11) & tmp12);
		when pcfar =>	pcnew := B & A;
		end case;

		------- reset overrides instruction fetch -----
		if reset='1' then
			romaddress <= "0000000000000000";
			pcnew := "0000000000000000";
		end if;
		
		romaddress <= pcnew;


		--------- synchronious stage (modify registers) -------
		if rising_edge(clk) then
			PC := pcnew;
			if reset='1' then
				SP := "11111111";
				O := (others => "11111111");
				R := "00000000";
				FETCHB := '0';
			else
				case SPCHANGE is
				when spnop  => 
				when spinc  => SP := SP + 1;
				when spdec  => SP := SP - 1; 
				when spdecx => SP := SP - x; 
				end case;
				if WRITEOUT then 
					O(x) := B;
				end if;
				R := R_NEW;
				FETCHB := FETCHB_NEW;
			end if;
		end if;

		

		
		----------------------- port output --------------		
		output <= O;

		--------------------- debug output --------------------
		test_pc <= PC;
		test_sp <= SP;
		test_r <= R;
		test_fetchb <= FETCHB;
	end process;
end rtl;
